module sprite_table(		input clk,

							output logic [0:15][0:15][0:3] enemy_0_0,
							output logic [0:15][0:15][0:3] enemy_0_1,
							output logic [0:15][0:15][0:3] enemy_1_0,
							output logic [0:15][0:15][0:3] enemy_1_1,
							output logic [0:15][0:15][0:3] enemy_2_0,
							output logic [0:15][0:15][0:3] enemy_2_1,
							output logic [0:15][0:15][0:3] enemy_3_0,
							output logic [0:15][0:15][0:3] enemy_3_1,
							output logic [0:15][0:15][0:3] enemy_4_00,
							output logic [0:15][0:15][0:3] enemy_5_00,
							output logic [0:15][0:15][0:3] enemy_6_00,
							output logic [0:15][0:15][0:3] enemy_7_00,
							output logic [0:15][0:15][0:3] enemy_8_0,
							output logic [0:15][0:15][0:3] enemy_8_1,
							output logic [0:15][0:15][0:3] enemy_8_2,
							output logic [0:15][0:15][0:3] enemy_9_00,
							output logic [0:15][0:15][0:3] player,
							output logic [0:15][0:15][0:3] player_missile,
							output logic [0:43][0:143][0:3] Logo_Galaxian,
							output logic [0:9][0:82][0:3] Logo_Gameover,
							output logic [0:8][0:119][0:3] Logo_Credits,
							output logic [0:8][0:136][0:3] Logo_Retry,
							output logic [0:31][0:31][0:3] explosion_0,
							output logic [0:31][0:31][0:3] explosion_1,
							output logic [0:31][0:31][0:3] explosion_2,
							output logic [0:31][0:31][0:3] explosion_3
					);	

	always_comb

	begin 

player <= 
'{ 
'{0,0,0,0,0,0,0,5,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,5,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,5,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,5,5,5,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,5,5,5,0,0,0,0,0,0,0},
'{0,0,0,6,0,0,5,5,5,0,0,6,0,0,0,0},
'{0,0,0,6,0,0,5,5,5,0,0,6,0,0,0,0},
'{0,0,0,5,0,5,5,5,5,5,0,5,0,0,0,0},
'{6,0,0,5,2,5,5,6,5,5,2,5,0,0,6,0},
'{6,0,0,2,5,5,6,6,6,5,5,2,0,0,6,0},
'{5,0,0,5,5,5,6,5,6,5,5,5,0,0,5,0},
'{5,0,5,5,5,5,5,5,5,5,5,5,5,0,5,0},
'{5,5,5,5,5,6,5,5,5,6,5,5,5,5,5,0},
'{5,5,5,0,6,6,5,5,5,6,6,0,5,5,5,0},
'{5,5,0,0,6,6,0,5,0,6,6,0,0,5,5,0},
'{5,0,0,0,0,0,0,5,0,0,0,0,0,0,5,0}
};

player_missile <= 
'{ 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 6, 6, 6, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 6, 3, 6, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 } 
};

enemy_0_0 <= 
'{ 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 6, 0, 0, 2, 0, 2, 0, 0, 6, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 6, 0, 5, 6, 5, 6, 5, 0, 6, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 6, 0, 5, 5, 5, 5, 5, 0, 6, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 6, 6, 6, 5, 5, 5, 6, 6, 6, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 6, 2, 2, 2, 6, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 6, 6, 6, 2, 2, 2, 6, 6, 6, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 6, 6, 6, 5, 5, 5, 6, 6, 6, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 6, 6, 0, 2, 2, 2, 0, 6, 6, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 6, 6, 0, 0, 2, 0, 0, 6, 6, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 } 
};

enemy_0_1 <= 
'{ 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 6, 0, 0, 2, 0, 2, 0, 0, 6, 0, 0, 0 }, 
'{ 0, 0, 6, 6, 6, 0, 0, 2, 0, 2, 0, 0, 6, 6, 6, 0 }, 
'{ 0, 0, 6, 6, 6, 0, 5, 6, 5, 6, 5, 0, 6, 6, 6, 0 }, 
'{ 0, 0, 6, 6, 6, 0, 5, 5, 5, 5, 5, 0, 6, 6, 6, 0 }, 
'{ 0, 0, 0, 6, 6, 6, 6, 5, 5, 5, 6, 6, 6, 6, 0, 0 }, 
'{ 0, 0, 0, 0, 6, 6, 6, 2, 2, 2, 6, 6, 6, 0, 0, 0 }, 
'{ 0, 0, 0, 6, 6, 6, 6, 2, 2, 2, 6, 6, 6, 6, 0, 0 }, 
'{ 0, 0, 6, 6, 6, 6, 6, 5, 5, 5, 6, 6, 6, 6, 6, 0 }, 
'{ 0, 0, 0, 6, 6, 6, 0, 2, 2, 2, 0, 6, 6, 6, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 } 
};

enemy_1_0 <= 
'{ 
'{ 0, 0, 0, 0, 0, 0, 13, 0, 13, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 13, 13, 10, 10, 13, 10, 10, 13, 13, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 13, 10, 10, 13, 10, 10, 13, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 13, 13, 13, 13, 13, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 13, 13, 11, 11, 13, 11, 11, 13, 13, 0, 0, 0, 0 }, 
'{ 0, 0, 13, 13, 13, 11, 11, 11, 11, 11, 13, 13, 13, 0, 0, 0 }, 
'{ 13, 13, 13, 13, 13, 11, 11, 11, 11, 11, 13, 13, 13, 13, 13, 0 }, 
'{ 0, 13, 13, 13, 0, 11, 11, 11, 11, 11, 0, 13, 13, 13, 0, 0 }, 
'{ 0, 0, 13, 13, 0, 0, 10, 0, 10, 0, 0, 13, 13, 0, 0, 0 }, 
'{ 0, 0, 13, 13, 0, 0, 10, 0, 10, 0, 0, 13, 13, 0, 0, 0 }, 
'{ 0, 0, 13, 13, 13, 0, 0, 0, 0, 0, 13, 13, 13, 0, 0, 0 }, 
'{ 0, 0, 0, 13, 13, 0, 0, 0, 0, 0, 13, 13, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 13, 13, 0, 0, 0, 13, 13, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 13, 13, 0, 13, 13, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 13, 0, 13, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 } 
};

enemy_1_1 <= 
'{ 
'{ 0, 0, 0, 0, 0, 0, 13, 0, 13, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 13, 0, 13, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 13, 13, 10, 10, 13, 10, 10, 13, 13, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 13, 10, 10, 13, 10, 10, 13, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 13, 13, 13, 13, 13, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 13, 11, 11, 13, 11, 11, 13, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 13, 13, 13, 11, 11, 11, 11, 11, 13, 13, 13, 0, 0, 0 }, 
'{ 13, 13, 13, 13, 13, 11, 11, 11, 11, 11, 13, 13, 13, 13, 13, 0 }, 
'{ 0, 13, 13, 13, 13, 11, 11, 11, 11, 11, 13, 13, 13, 13, 0, 0 }, 
'{ 0, 13, 10, 13, 13, 0, 10, 0, 10, 0, 13, 13, 10, 13, 0, 0 }, 
'{ 13, 13, 10, 13, 0, 0, 10, 0, 10, 0, 0, 13, 10, 13, 13, 0 }, 
'{ 13, 10, 13, 13, 0, 0, 0, 0, 0, 0, 0, 13, 13, 10, 13, 0 }, 
'{ 13, 10, 10, 13, 0, 0, 0, 0, 0, 0, 0, 13, 10, 10, 13, 0 }, 
'{ 13, 10, 10, 13, 0, 0, 0, 0, 0, 0, 0, 13, 10, 10, 13, 0 }, 
'{ 13, 13, 13, 13, 0, 0, 0, 0, 0, 0, 0, 13, 13, 13, 13, 0 }, 
'{ 0, 13, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 13, 0, 0 } 
};

enemy_2_0 <= 
'{ 
'{ 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 1, 1, 8, 8, 1, 8, 8, 1, 1, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 1, 8, 8, 1, 8, 8, 1, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 1, 1, 12, 12, 1, 12, 12, 1, 1, 0, 0, 0, 0 }, 
'{ 0, 0, 1, 1, 1, 12, 12, 12, 12, 12, 1, 1, 1, 0, 0, 0 }, 
'{ 1, 1, 1, 1, 1, 12, 12, 12, 12, 12, 1, 1, 1, 1, 1, 0 }, 
'{ 0, 1, 1, 1, 0, 12, 12, 12, 12, 12, 0, 1, 1, 1, 0, 0 }, 
'{ 0, 0, 1, 1, 0, 0, 8, 0, 8, 0, 0, 1, 1, 0, 0, 0 }, 
'{ 0, 0, 1, 1, 0, 0, 8, 0, 8, 0, 0, 1, 1, 0, 0, 0 }, 
'{ 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0 }, 
'{ 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 } 
};

enemy_2_1 <= 
'{ 
'{ 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 1, 1, 8, 8, 1, 8, 8, 1, 1, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 1, 8, 8, 1, 8, 8, 1, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 1, 12, 12, 1, 12, 12, 1, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 1, 1, 1, 12, 12, 12, 12, 12, 1, 1, 1, 0, 0, 0 }, 
'{ 1, 1, 1, 1, 1, 12, 12, 12, 12, 12, 1, 1, 1, 1, 1, 0 }, 
'{ 0, 1, 1, 1, 1, 12, 12, 12, 12, 12, 1, 1, 1, 1, 0, 0 }, 
'{ 0, 1, 8, 1, 1, 0, 8, 0, 8, 0, 1, 1, 8, 1, 0, 0 }, 
'{ 1, 1, 8, 1, 0, 0, 8, 0, 8, 0, 0, 1, 8, 1, 1, 0 }, 
'{ 1, 8, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 8, 1, 0 }, 
'{ 1, 8, 8, 1, 0, 0, 0, 0, 0, 0, 0, 1, 8, 8, 1, 0 }, 
'{ 1, 8, 8, 1, 0, 0, 0, 0, 0, 0, 0, 1, 8, 8, 1, 0 }, 
'{ 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0 }, 
'{ 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0 } 
};

enemy_3_0 <= 
'{ 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 1, 0, 0, 0, 11, 0, 0, 0, 1, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 1, 0, 11, 6, 11, 6, 11, 0, 1, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 1, 6, 6, 11, 6, 6, 1, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 11, 11, 11, 11, 11, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 1, 1, 11, 11, 11, 1, 1, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 1, 1, 6, 6, 6, 1, 1, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 1, 1, 0, 6, 6, 6, 0, 1, 1, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 1, 1, 0, 11, 11, 11, 0, 1, 1, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 1, 1, 0, 6, 6, 6, 0, 1, 1, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 1, 1, 0, 0, 6, 0, 0, 1, 1, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 } 
};

enemy_3_1 <= 
'{ 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 1, 0, 0, 0, 0, 11, 0, 0, 0, 0, 1, 0, 0, 0 }, 
'{ 0, 0, 0, 1, 0, 11, 6, 11, 6, 11, 0, 1, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 1, 6, 6, 11, 6, 6, 1, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 11, 11, 11, 11, 11, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 1, 1, 11, 11, 11, 1, 1, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 1, 1, 1, 6, 6, 6, 1, 1, 1, 0, 0, 0, 0 }, 
'{ 0, 0, 1, 1, 1, 0, 6, 6, 6, 0, 1, 1, 1, 0, 0, 0 }, 
'{ 0, 1, 1, 1, 1, 0, 11, 11, 11, 0, 1, 1, 1, 1, 0, 0 }, 
'{ 0, 1, 1, 1, 0, 0, 6, 6, 6, 0, 0, 1, 1, 1, 0, 0 }, 
'{ 0, 1, 1, 1, 0, 0, 0, 6, 0, 0, 0, 1, 1, 1, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 } 
};

enemy_4_00 <= 
'{ 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 1, 0, 0, 0, 10, 10, 10, 0, 0, 0, 1, 0, 0, 0 }, 
'{ 0, 0, 1, 0, 0, 10, 10, 10, 10, 10, 0, 0, 1, 0, 0, 0 }, 
'{ 0, 0, 1, 11, 10, 10, 11, 10, 11, 10, 10, 11, 1, 0, 0, 0 }, 
'{ 0, 0, 1, 11, 11, 11, 11, 10, 11, 11, 11, 11, 1, 0, 0, 0 }, 
'{ 0, 0, 1, 1, 11, 11, 11, 11, 11, 11, 11, 1, 1, 0, 0, 0 }, 
'{ 0, 0, 0, 1, 1, 11, 0, 11, 0, 11, 1, 1, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 1, 1, 0, 11, 0, 1, 1, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 1, 0, 11, 0, 1, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 } 
};

enemy_5_00 <= 
'{ 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 6, 0, 6, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 3, 0, 3, 0, 6, 0, 6, 0, 3, 0, 3, 0, 0, 0 }, 
'{ 0, 0, 3, 3, 3, 0, 0, 9, 0, 0, 3, 3, 3, 0, 0, 0 }, 
'{ 0, 0, 0, 3, 3, 0, 9, 9, 9, 0, 3, 3, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 3, 3, 0, 9, 9, 9, 0, 3, 3, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 3, 3, 9, 9, 9, 3, 3, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 9, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 9, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 } 
};

enemy_6_00 <= 
'{ 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 8, 8, 7, 8, 8, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 8, 8, 7, 7, 7, 8, 8, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 8, 7, 7, 6, 7, 7, 8, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 7, 7, 7, 7, 6, 7, 7, 7, 7, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 7, 7, 7, 6, 6, 6, 7, 7, 7, 0, 0, 0, 0 }, 
'{ 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0 }, 
'{ 0, 0, 7, 7, 0, 0, 7, 7, 7, 0, 0, 7, 7, 0, 0, 0 }, 
'{ 0, 0, 7, 0, 0, 0, 0, 7, 0, 0, 0, 0, 7, 0, 0, 0 }, 
'{ 0, 0, 7, 0, 0, 0, 0, 7, 0, 0, 0, 0, 7, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 } 
};

enemy_7_00 <= 
'{ 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 6, 6, 0, 6, 6, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 6, 1, 6, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 1, 1, 1, 1, 1, 1, 0, 1, 0, 1, 1, 1, 1, 1, 1, 0 }, 
'{ 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0 }, 
'{ 0, 5, 5, 5, 5, 5, 5, 1, 5, 5, 5, 5, 5, 5, 0, 0 }, 
'{ 0, 0, 0, 5, 5, 5, 0, 1, 0, 5, 5, 5, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 } 
};

enemy_8_0 <= 
'{ 
'{ 0, 0, 0, 0, 0, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 6, 6, 0, 0, 0, 0, 1, 5, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 6, 6, 6, 0, 0, 1, 5, 5, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 6, 6, 6, 1, 1, 5, 5, 0, 0, 0 }, 
'{ 0, 6, 6, 6, 6, 0, 0, 6, 1, 1, 5, 5, 5, 0, 0, 0 }, 
'{ 0, 0, 6, 6, 6, 6, 6, 1, 1, 1, 5, 5, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 6, 6, 6, 6, 6, 1, 5, 5, 5, 6, 6, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 6, 6, 5, 5, 5, 5, 6, 6, 6, 6 }, 
'{ 0, 0, 0, 0, 0, 0, 1, 5, 6, 6, 6, 0, 0, 6, 6, 6 }, 
'{ 0, 0, 0, 0, 0, 0, 1, 5, 5, 6, 6, 6, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 1, 0, 0, 0, 6, 6, 6, 0, 0, 0, 0 }, 
'{ 0, 0, 1, 0, 1, 0, 0, 0, 0, 6, 6, 6, 6, 0, 0, 0 }, 
'{ 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 6, 6, 6, 0, 0, 0 }, 
'{ 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 6, 6, 6, 6, 0, 0 }, 
'{ 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 } 
};

enemy_8_1 <= 
'{ 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 6, 6, 6, 0, 0, 0, 0, 0, 0, 1, 5, 0, 0, 0 }, 
'{ 0, 0, 0, 6, 6, 6, 6, 0, 0, 0, 1, 5, 5, 6, 0, 0 }, 
'{ 0, 0, 0, 0, 6, 6, 6, 6, 0, 1, 1, 5, 6, 6, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 6, 6, 6, 1, 1, 5, 5, 6, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 5, 5, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 6, 6, 1, 1, 5, 6, 6, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 6, 6, 6, 6, 5, 6, 6, 6, 6, 0, 0 }, 
'{ 0, 0, 0, 0, 6, 6, 6, 6, 6, 5, 0, 6, 6, 6, 6, 0 }, 
'{ 0, 0, 0, 6, 6, 6, 6, 6, 0, 0, 0, 0, 6, 6, 6, 6 }, 
'{ 0, 0, 0, 6, 6, 6, 6, 0, 0, 0, 0, 0, 0, 6, 6, 0 }, 
'{ 0, 1, 0, 6, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 } 
};

enemy_8_2 <= 
'{ 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 1, 5, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 1, 5, 5, 0, 0, 0 }, 
'{ 6, 6, 6, 6, 6, 0, 0, 0, 6, 1, 5, 5, 0, 0, 0, 0 }, 
'{ 0, 6, 6, 6, 6, 6, 6, 0, 1, 1, 5, 5, 0, 0, 0, 0 }, 
'{ 0, 0, 6, 6, 6, 6, 6, 1, 1, 5, 5, 5, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 6, 6, 6, 1, 5, 5, 5, 6, 6, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 1, 1, 5, 5, 5, 6, 6, 6, 6, 0 }, 
'{ 0, 0, 0, 0, 0, 1, 5, 6, 6, 6, 5, 6, 6, 6, 6, 6 }, 
'{ 0, 0, 0, 0, 0, 1, 6, 6, 6, 6, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 1, 0, 6, 6, 6, 6, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 1, 0, 1, 0, 0, 6, 6, 6, 6, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 1, 0, 0, 0, 6, 6, 6, 6, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 1, 0, 1, 0, 0, 6, 6, 6, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 1, 0, 0, 0, 0, 0, 0, 6, 6, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 } 
};

enemy_9_00 <= 
'{ 
'{ 0, 0, 0, 0, 0, 1, 1, 5, 1, 1, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 1, 1, 1, 5, 1, 1, 1, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 1, 1, 1, 1, 5, 1, 1, 1, 1, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 1, 1, 1, 6, 6, 6, 1, 1, 1, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 1, 1, 6, 6, 5, 6, 6, 1, 1, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 1, 1, 1, 6, 6, 6, 1, 1, 1, 0, 0, 0, 0 }, 
'{ 0, 5, 0, 1, 1, 1, 1, 6, 1, 1, 1, 1, 0, 5, 0, 0 }, 
'{ 0, 1, 1, 0, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 0, 0 }, 
'{ 0, 1, 1, 0, 0, 1, 1, 6, 1, 1, 0, 0, 1, 1, 0, 0 }, 
'{ 0, 1, 1, 6, 0, 0, 0, 6, 0, 0, 0, 6, 1, 1, 0, 0 }, 
'{ 0, 1, 1, 6, 6, 0, 1, 6, 1, 0, 6, 6, 1, 1, 0, 0 }, 
'{ 0, 1, 1, 6, 6, 6, 1, 6, 1, 6, 6, 6, 1, 1, 0, 0 }, 
'{ 0, 1, 1, 0, 6, 6, 1, 1, 1, 6, 6, 0, 1, 1, 0, 0 }, 
'{ 0, 1, 1, 0, 0, 6, 1, 1, 1, 6, 0, 0, 1, 1, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 5, 1, 5, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 5, 1, 5, 0, 0, 0, 0, 0, 0, 0 } 
};



Logo_Galaxian <= 
'{ 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 9, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 9, 9, 9, 9, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 9, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 9, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 9, 9, 9, 9, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 9, 9, 9, 0, 0, 0, 0, 0, 9, 9, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 9, 0, 0, 0, 0, 0, 0, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 9, 9, 9, 9, 2, 2, 2, 2, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 9, 9, 0, 0, 0, 0, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 9, 2, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 9, 2, 2, 2, 2, 2, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 0, 0, 0, 0, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 9, 0, 0, 0, 0, 9, 9, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 9, 9, 2, 2, 2, 2, 2, 9, 9, 9, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 0, 0, 0, 9, 9, 9, 2, 2, 2, 2, 2, 9, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 0, 0, 0, 0, 0, 0, 0, 9, 9, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 0, 0, 0, 9, 2, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 0, 0, 0, 0, 0, 0, 9, 9, 9, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 9, 9, 2, 9, 9, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 0, 0, 0, 0, 0, 0, 9, 9, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 0, 0, 0, 0, 9, 9, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 9, 0, 0, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 0, 0, 0, 9, 9, 2, 2, 2, 2, 9, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 0, 0, 0, 9, 2, 2, 9, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 2, 2, 2, 2, 2, 2, 9, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 0, 0, 9, 9, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 9, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 0, 0, 0, 0, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 9, 2, 2, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 2, 2, 2, 2, 9, 0, 0, 0, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 9, 9, 9, 9, 2, 2, 2, 2, 2, 9, 0, 0, 9, 2, 2, 2, 2, 2, 2, 9, 9, 0, 0, 0, 0, 0, 9, 9, 9, 9, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 9, 9, 9, 9, 9, 0, 0, 0, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 9, 9, 9, 9, 9, 9, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2, 9, 9, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 9, 9, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 9, 2, 2, 2, 9, 9, 9, 9, 0, 0, 0, 0, 0, 9, 9, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 9, 0, 0, 0, 0, 9, 9, 9, 9, 9, 9, 2, 2, 2, 2, 2, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 9, 9, 9, 9, 9, 9, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 9, 9, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 9, 9, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 9, 0, 0, 0, 0, 0, 9, 2, 9, 9, 0, 0, 0, 0, 0, 9, 9, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 2, 2, 2, 2, 2, 2, 9, 9, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 9, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 9, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 9, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 9, 0, 0, 0, 0, 0, 0, 9, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 9, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 9, 0, 0, 0, 0, 0, 0, 9, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 9, 0, 0, 0, 0, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 9, 2, 9, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 9, 9, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 9, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 9, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 9, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 2, 9, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 9, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 0, 0, 0, 0, 9, 9, 9, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 9, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 9, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 9, 9, 9, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 9, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 0, 0, 9, 9, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 9, 2, 2, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 0, 0, 9, 9, 9, 9, 2, 2, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 2, 2, 2, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 2, 2, 9, 9, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 9, 9, 9, 9, 0, 0, 9, 9, 9, 9, 2, 2, 2, 2, 9, 9, 0, 0, 0, 0, 0, 0, 0, 9, 9, 9, 9, 0, 0, 9, 9, 9, 0, 0, 0, 0, 0, 9, 2, 9, 9, 9, 0, 0, 0, 0, 0, 0, 9, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 9, 9, 9, 9, 9, 9, 9, 2, 2, 2, 2, 9, 9, 2, 2, 2, 9, 9, 9, 9, 9, 2, 2, 2, 2, 2, 9, 9, 9, 9, 9, 9, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 }, 
'{ 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 } 
};
 
Logo_Gameover <= 
'{ 
'{ 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 0, 7, 7, 7, 0, 0, 0, 0, 7, 7, 7, 0, 0, 0, 7, 7, 7, 0, 0, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 0, 0, 0, 7, 7, 0, 0, 0, 7, 7, 0, 0, 7, 7, 7, 7, 7, 7, 7, 0, 0, 7, 7, 7, 7, 7, 7, 7, 0, 0, 7, 7, 0 }, 
'{ 7, 7, 7, 0, 0, 7, 7, 7, 0, 0, 0, 0, 7, 7, 7, 7, 0, 0, 0, 7, 7, 7, 0, 0, 0, 7, 7, 7, 0, 0, 7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 7, 0, 0, 0, 7, 7, 0, 0, 7, 7, 0, 0, 0, 7, 7, 0, 0, 7, 7, 0, 0, 0, 0, 0, 0, 0, 7, 7, 0, 0, 0, 7, 7, 7, 0, 7, 7, 0 }, 
'{ 7, 7, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 7, 7, 7, 7, 0, 0, 0, 7, 7, 7, 0, 0, 0, 7, 7, 7, 0, 0, 7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 0, 0, 0, 0, 7, 7, 0, 0, 7, 7, 0, 0, 0, 7, 7, 0, 0, 7, 7, 0, 0, 0, 0, 0, 0, 0, 7, 7, 0, 0, 0, 0, 7, 7, 0, 7, 7, 0 }, 
'{ 7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 0, 7, 7, 0, 0, 0, 7, 7, 7, 7, 0, 7, 7, 7, 7, 0, 0, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 0, 0, 0, 7, 7, 0, 0, 0, 0, 7, 7, 0, 0, 0, 7, 0, 0, 7, 7, 0, 0, 0, 7, 7, 7, 7, 7, 7, 0, 0, 0, 7, 7, 0, 0, 0, 7, 7, 0, 0, 0, 7, 0 }, 
'{ 7, 7, 0, 0, 7, 7, 7, 7, 0, 0, 0, 7, 7, 0, 0, 7, 7, 0, 0, 7, 7, 0, 7, 0, 7, 0, 7, 7, 0, 0, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 0, 0, 0, 7, 7, 0, 0, 0, 0, 0, 7, 7, 0, 0, 7, 7, 0, 7, 7, 0, 0, 0, 7, 7, 7, 7, 7, 7, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 7, 0 }, 
'{ 7, 7, 0, 0, 0, 7, 7, 7, 0, 0, 0, 7, 7, 7, 7, 7, 7, 0, 0, 7, 7, 0, 7, 0, 7, 0, 7, 7, 0, 0, 7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 0, 0, 0, 0, 7, 7, 0, 0, 0, 7, 7, 0, 7, 0, 0, 0, 0, 7, 7, 0, 0, 0, 0, 0, 0, 0, 7, 7, 0, 0, 0, 7, 7, 0, 0, 0, 7, 0 }, 
'{ 7, 7, 0, 0, 0, 0, 7, 7, 0, 0, 7, 7, 7, 7, 7, 7, 7, 0, 0, 7, 7, 0, 7, 7, 7, 0, 7, 7, 0, 0, 7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 0, 0, 0, 0, 7, 7, 0, 0, 0, 0, 7, 7, 7, 0, 0, 0, 0, 7, 7, 0, 0, 0, 0, 0, 0, 0, 7, 7, 0, 0, 0, 7, 7, 0, 0, 0, 0, 0 }, 
'{ 0, 7, 7, 7, 7, 7, 7, 7, 0, 0, 7, 7, 0, 0, 0, 0, 7, 7, 0, 7, 7, 0, 7, 7, 7, 0, 7, 7, 0, 0, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 0, 0, 0, 7, 7, 7, 0, 7, 7, 7, 0, 0, 0, 0, 7, 7, 7, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 0, 0, 7, 7, 0, 0, 0, 7, 7, 0, 0, 0, 7, 0 }, 
'{ 0, 0, 7, 7, 7, 7, 0, 7, 0, 0, 7, 7, 0, 0, 0, 0, 7, 7, 0, 7, 7, 0, 7, 7, 7, 0, 7, 7, 0, 0, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7, 0, 0, 0, 0, 0, 7, 7, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 0, 0, 7, 7, 0, 0, 0, 0, 7, 7, 0, 7, 7, 0 } 
};

Logo_Retry <= 
'{ 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 11, 10, 10, 9, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 11, 0, 0, 10, 10, 0, 10, 9, 9, 9, 10, 0, 10, 10, 10, 9, 0, 0, 9, 10, 10, 10, 0, 0, 9, 10, 10, 10, 0, 0, 0, 0, 0, 0, 0, 9, 0, 10, 10, 0, 9, 0, 0, 0, 0, 0, 0, 0, 10, 11, 10, 10, 0, 0, 9, 10, 10, 9, 0, 0, 0, 0, 0, 0, 0, 0, 10, 11, 10, 10, 0, 0, 10, 9, 9, 9, 10, 0, 9, 0, 0, 10, 10, 0, 0, 0, 0, 0, 0, 0, 10, 10, 10, 9, 0, 0, 9, 10, 10, 11, 0, 0, 10, 10, 10, 9, 0, 0, 10, 10, 9, 0, 0, 0, 11, 9, 10, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 11, 0, 0, 9, 0, 0, 10, 10, 0, 0, 0, 0, 9, 0, 0, 9, 0, 0, 9, 10, 0, 0, 0, 0, 9, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 9, 9, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 9, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 10, 10, 0, 0, 0, 0, 9, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 9, 0, 0, 9, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 9, 0, 0, 0, 11, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 11, 9, 10, 0, 0, 0, 10, 10, 0, 0, 0, 0, 11, 10, 10, 10, 0, 0, 0, 10, 9, 10, 0, 0, 0, 10, 9, 10, 0, 0, 0, 0, 0, 0, 0, 0, 10, 9, 9, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 10, 10, 0, 0, 10, 10, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 10, 10, 0, 0, 0, 0, 0, 9, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 10, 10, 10, 11, 0, 0, 9, 0, 0, 9, 0, 0, 10, 10, 10, 11, 0, 0, 0, 0, 9, 0, 0, 0, 9, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 11, 0, 0, 0, 0, 0, 10, 10, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 9, 10, 10, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 9, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 10, 10, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 11, 0, 0, 11, 0, 0, 11, 0, 0, 9, 0, 0, 11, 0, 0, 0, 0, 9, 0, 0, 0, 9, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 11, 0, 0, 0, 0, 0, 10, 10, 0, 0, 0, 0, 0, 9, 9, 9, 0, 0, 9, 9, 9, 10, 0, 0, 9, 9, 9, 10, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 9, 9, 0, 0, 10, 9, 9, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 9, 9, 0, 0, 10, 10, 0, 0, 0, 0, 0, 10, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 10, 9, 10, 0, 10, 9, 9, 9, 0, 0, 9, 9, 10, 9, 10, 0, 0, 0, 9, 0, 0, 0, 9, 0, 0, 9, 0, 0, 0, 9, 9, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 9, 9, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 9, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 } 
};

Logo_Credits <= 
'{ 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 9, 9, 10, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0 }, 
'{ 0, 0, 11, 10, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 10, 0, 0, 0, 11, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 10, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 10, 10, 0, 0, 0, 0, 0, 0, 0, 0, 10, 9, 0, 0, 9, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0 }, 
'{ 0, 0, 9, 0, 0, 11, 0, 0, 9, 0, 0, 10, 10, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 10, 0, 0, 10, 11, 10, 10, 0, 0, 11, 0, 10, 10, 0, 0, 10, 10, 10, 9, 0, 0, 10, 9, 9, 9, 10, 0, 9, 10, 10, 10, 0, 0, 11, 9, 11, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 10, 0, 0, 0, 0, 0, 0, 0, 0, 10, 9, 0, 0, 9, 10, 0, 10, 10, 9, 0, 0, 0, 10, 9, 10, 10, 0, 0, 11, 9, 10, 11, 0, 0, 10, 10, 10, 9, 0, 0, 10, 10, 10, 9, 0, 0, 0, 0, 9, 0 }, 
'{ 0, 0, 11, 10, 9, 0, 0, 0, 9, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 10, 0, 0, 0, 11, 0, 0, 0, 0, 11, 10, 9, 0, 0, 0, 0, 0, 0, 9, 0, 0, 10, 10, 0, 0, 0, 0, 9, 10, 0, 0, 0, 0, 11, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 0, 0, 9, 0, 0, 0, 0, 0, 0, 10, 0, 10, 10, 0, 10, 0, 0, 0, 9, 0, 0, 0, 9, 0, 0, 0, 0, 0, 11, 0, 0, 9, 0, 0, 0, 0, 0, 9, 0, 0, 9, 0, 0, 9, 0, 0, 0, 0, 9, 0 }, 
'{ 0, 0, 9, 0, 0, 9, 0, 0, 0, 9, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 10, 0, 0, 0, 11, 0, 0, 0, 0, 11, 9, 10, 0, 0, 0, 10, 10, 10, 11, 0, 0, 10, 10, 0, 0, 0, 0, 0, 10, 9, 10, 0, 0, 9, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 11, 0, 9, 0, 0, 0, 0, 0, 0, 10, 0, 9, 9, 0, 10, 0, 0, 0, 9, 0, 0, 0, 11, 0, 0, 0, 0, 0, 9, 0, 0, 9, 0, 0, 10, 10, 10, 11, 0, 0, 11, 10, 10, 10, 0, 0, 0, 0, 9, 0 }, 
'{ 0, 0, 9, 0, 0, 9, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 9, 0, 0, 0, 9, 0, 0, 0, 0, 11, 0, 9, 10, 0, 0, 9, 0, 0, 11, 0, 0, 10, 10, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 9, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 9, 10, 0, 10, 11, 0, 0, 0, 0, 0, 0, 0, 10, 0, 10, 0, 0, 10, 0, 0, 0, 9, 0, 0, 0, 9, 0, 0, 0, 0, 0, 9, 0, 0, 9, 0, 0, 9, 0, 0, 11, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 9, 0 }, 
'{ 0, 0, 11, 9, 9, 9, 0, 0, 0, 10, 10, 0, 0, 0, 0, 0, 0, 0, 0, 7, 10, 9, 9, 10, 0, 0, 0, 10, 9, 9, 0, 0, 11, 0, 0, 9, 0, 0, 9, 9, 10, 9, 10, 0, 10, 10, 0, 0, 0, 0, 9, 9, 9, 10, 0, 0, 9, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 9, 9, 10, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 10, 0, 0, 0, 9, 0, 0, 0, 0, 9, 9, 9, 0, 0, 9, 0, 0, 9, 0, 0, 9, 9, 10, 9, 10, 0, 0, 9, 9, 9, 0, 0, 0, 0, 9, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 } 
};

explosion_0 <= 
'{ 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 3, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 3, 3, 0, 3, 3, 5, 5, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 5, 5, 0, 0, 3, 0, 3, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 3, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 5, 3, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 3, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 3, 6, 0, 3, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 3, 0, 0, 3, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 3, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 3, 5, 0, 5, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 6, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 3, 0, 3, 5, 0, 0, 0, 0, 0, 6, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 6, 6, 6, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 3, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 6, 0, 0, 6, 6, 6, 0, 0, 6, 0, 0, 0, 0, 0, 3, 0, 0, 3, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 6, 0, 0, 6, 6, 6, 0, 0, 6, 0, 0, 0, 0, 0, 3, 0, 5, 0, 3, 0, 0, 0 }, 
'{ 0, 0, 0, 3, 0, 6, 0, 0, 0, 0, 6, 0, 6, 6, 6, 6, 6, 0, 6, 0, 0, 0, 0, 0, 6, 3, 0, 0, 3, 0, 0, 0 }, 
'{ 0, 0, 3, 0, 3, 0, 0, 6, 0, 0, 6, 0, 6, 6, 6, 6, 6, 0, 6, 0, 0, 6, 0, 0, 0, 3, 0, 3, 0, 0, 0, 0 }, 
'{ 0, 0, 3, 0, 3, 0, 0, 6, 0, 0, 6, 6, 6, 6, 6, 6, 6, 6, 6, 0, 0, 6, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0 }, 
'{ 0, 5, 5, 5, 5, 0, 0, 6, 0, 0, 6, 6, 6, 6, 6, 6, 6, 6, 6, 0, 0, 6, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0 }, 
'{ 3, 0, 0, 0, 0, 0, 0, 6, 0, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 0, 6, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0 }, 
'{ 3, 0, 0, 0, 3, 0, 0, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0 }, 
'{ 0, 5, 5, 5, 3, 0, 0, 6, 6, 6, 0, 6, 6, 6, 6, 6, 6, 6, 0, 6, 6, 6, 0, 0, 5, 0, 5, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 3, 3, 3, 6, 0, 6, 6, 0, 0, 6, 6, 0, 6, 0, 6, 6, 0, 0, 6, 6, 0, 0, 5, 0, 0, 3, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 3, 3, 0, 3, 6, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 6, 0, 6, 0, 3, 0, 3, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 3, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 3, 3, 0, 0, 3, 0, 0, 0, 0, 0, 3, 0, 0, 3, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 3, 0, 0, 6, 0, 0, 0, 0, 6, 0, 0, 3, 0, 0, 6, 6, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 5, 0, 0, 0, 3, 0, 0, 5, 5, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 3, 3, 3, 3, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 } 
};

explosion_1 <= 
'{ 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0 }, 
'{ 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 3, 3, 3, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 3, 3, 0, 0, 0, 0, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 6, 0, 0, 0, 3, 3, 3, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 3, 0, 6, 0, 0, 3, 3, 3, 3, 0, 6, 0, 3, 3, 0, 0, 0, 3, 3, 0, 3, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 3, 0, 0, 3, 3, 0, 6, 0, 3, 0, 3, 3, 3, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 3, 3, 0, 0, 0, 3, 3, 5, 0, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 5, 5, 5, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 3, 0, 3, 3, 3, 3, 3, 0, 3, 3, 0, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 6, 0, 0, 0, 3, 3, 3, 0, 3, 3, 3, 5, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 3, 3, 0, 0, 3, 3, 3, 3, 3, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 6, 3, 0, 3, 3, 0, 0, 3, 3, 3, 0, 0, 0 }, 
'{ 0, 0, 0, 3, 3, 3, 0, 3, 0, 5, 5, 0, 0, 5, 5, 5, 5, 0, 5, 3, 6, 3, 0, 3, 3, 0, 0, 3, 0, 0, 0, 0 }, 
'{ 0, 0, 3, 3, 3, 0, 3, 3, 5, 0, 5, 0, 5, 0, 5, 0, 0, 5, 5, 3, 3, 3, 0, 3, 3, 0, 0, 3, 3, 0, 0, 0 }, 
'{ 0, 0, 3, 3, 0, 3, 3, 3, 5, 5, 5, 5, 0, 5, 0, 5, 0, 5, 5, 5, 3, 0, 3, 3, 3, 0, 5, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 3, 3, 0, 3, 3, 3, 0, 5, 5, 3, 0, 0, 6, 5, 0, 0, 0, 5, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 3, 3, 0, 3, 3, 3, 0, 0, 0, 0, 5, 5, 5, 5, 5, 5, 0, 0, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 3, 3, 0, 3, 3, 6, 5, 5, 5, 5, 0, 5, 6, 5, 0, 0, 0, 0, 5, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 3, 3, 3, 0, 3, 6, 5, 5, 5, 0, 0, 0, 5, 5, 6, 0, 5, 5, 5, 3, 0, 3, 3, 3, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 3, 3, 3, 3, 3, 5, 5, 0, 5, 5, 0, 5, 0, 5, 0, 5, 5, 5, 5, 3, 3, 0, 3, 3, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 3, 3, 3, 3, 0, 3, 5, 5, 0, 5, 0, 0, 0, 0, 0, 5, 5, 6, 5, 0, 3, 3, 3, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 3, 3, 3, 3, 0, 3, 5, 0, 0, 0, 5, 5, 0, 5, 5, 0, 5, 5, 5, 3, 0, 3, 3, 0, 6, 0, 0, 0, 0 }, 
'{ 0, 3, 0, 0, 3, 3, 0, 3, 3, 5, 0, 5, 5, 5, 5, 0, 5, 5, 5, 5, 3, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 3, 0, 0, 0, 3, 3, 3, 3, 3, 5, 6, 5, 3, 3, 3, 5, 6, 5, 3, 0, 3, 3, 3, 0, 3, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 3, 3, 0, 0, 3, 3, 0, 3, 3, 0, 3, 3, 3, 3, 0, 3, 3, 3, 0, 0, 5, 5, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 3, 0, 0, 5, 0, 0, 3, 3, 0, 0, 3, 3, 0, 3, 3, 3, 0, 3, 3, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 6, 0, 3, 0, 0, 3, 3, 3, 3, 3, 3, 0, 3, 3, 3, 3, 3, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 6, 0, 0, 3, 0, 0, 0, 3, 3, 0, 3, 3, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0 }, 
'{ 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 } 
};

explosion_2 <= 
'{ 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 3, 3, 3, 3, 3, 0, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 3 }, 
'{ 0, 3, 0, 0, 0, 0, 0, 0, 3, 3, 3, 3, 3, 3, 0, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 3, 0 }, 
'{ 0, 0, 3, 0, 0, 0, 0, 3, 3, 3, 3, 3, 3, 3, 0, 3, 3, 3, 3, 3, 0, 3, 0, 5, 5, 3, 3, 0, 3, 3, 0, 0 }, 
'{ 0, 0, 3, 3, 3, 0, 3, 3, 5, 5, 0, 0, 3, 3, 3, 3, 3, 5, 5, 0, 5, 0, 5, 0, 5, 5, 3, 0, 0, 0, 6, 0 }, 
'{ 0, 0, 0, 6, 0, 0, 3, 3, 5, 0, 5, 5, 0, 3, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 0, 5, 3, 3, 0, 6, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 5, 6, 5, 5, 5, 5, 0, 5, 5, 3, 5, 5, 5, 5, 3, 5, 5, 5, 0, 3, 3, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 3, 3, 5, 5, 5, 5, 5, 3, 5, 5, 5, 6, 6, 5, 5, 5, 5, 5, 3, 5, 5, 5, 0, 3, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 3, 5, 5, 0, 5, 3, 5, 5, 5, 3, 3, 3, 3, 5, 0, 5, 5, 5, 5, 5, 6, 5, 5, 0, 3, 3, 3, 0, 0 }, 
'{ 0, 0, 3, 3, 5, 0, 5, 5, 3, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 3, 5, 5, 6, 3, 5, 0, 5, 5, 5, 3, 3, 0 }, 
'{ 0, 3, 3, 5, 0, 5, 5, 3, 5, 5, 5, 5, 5, 0, 5, 5, 5, 0, 5, 5, 5, 5, 5, 3, 5, 5, 5, 5, 0, 3, 3, 0 }, 
'{ 0, 3, 3, 0, 5, 5, 5, 3, 5, 5, 0, 5, 5, 5, 0, 5, 5, 0, 5, 5, 5, 0, 5, 5, 5, 5, 3, 5, 3, 0, 3, 3 }, 
'{ 0, 3, 3, 0, 5, 5, 5, 5, 5, 5, 5, 0, 5, 6, 5, 5, 0, 5, 5, 5, 0, 5, 5, 0, 5, 5, 3, 5, 0, 3, 3, 0 }, 
'{ 0, 3, 3, 5, 0, 5, 6, 5, 5, 0, 0, 5, 0, 5, 0, 0, 0, 5, 0, 0, 0, 5, 3, 5, 0, 5, 3, 5, 5, 0, 3, 3 }, 
'{ 0, 0, 3, 5, 5, 3, 5, 5, 3, 5, 0, 0, 5, 0, 0, 5, 0, 0, 5, 0, 5, 5, 5, 5, 0, 5, 5, 5, 5, 0, 3, 3 }, 
'{ 0, 0, 3, 3, 5, 3, 5, 5, 3, 5, 5, 0, 0, 5, 0, 5, 0, 5, 0, 0, 5, 5, 5, 0, 5, 5, 5, 5, 0, 3, 3, 3 }, 
'{ 0, 0, 0, 3, 0, 5, 3, 5, 3, 5, 3, 0, 0, 0, 5, 5, 5, 5, 0, 0, 0, 5, 5, 5, 5, 5, 5, 0, 3, 3, 3, 0 }, 
'{ 0, 0, 3, 0, 3, 5, 5, 5, 5, 5, 0, 5, 6, 5, 5, 5, 5, 6, 5, 5, 0, 5, 5, 5, 6, 5, 0, 3, 3, 3, 0, 0 }, 
'{ 0, 0, 3, 3, 5, 6, 5, 5, 5, 0, 0, 0, 5, 0, 0, 5, 5, 0, 0, 0, 0, 0, 5, 5, 5, 5, 3, 3, 3, 0, 0, 0 }, 
'{ 0, 0, 3, 3, 5, 5, 3, 5, 5, 5, 5, 5, 0, 5, 0, 0, 5, 5, 0, 0, 5, 5, 5, 5, 5, 5, 3, 3, 0, 3, 0, 0 }, 
'{ 0, 0, 3, 3, 0, 5, 5, 3, 5, 5, 5, 0, 0, 5, 0, 0, 0, 5, 0, 5, 5, 5, 3, 5, 5, 6, 3, 3, 0, 3, 3, 0 }, 
'{ 0, 0, 0, 3, 3, 5, 5, 5, 5, 5, 5, 0, 5, 0, 0, 0, 0, 0, 0, 0, 5, 5, 5, 5, 5, 5, 3, 3, 0, 3, 0, 6 }, 
'{ 0, 0, 0, 0, 3, 0, 5, 5, 3, 5, 0, 0, 0, 5, 5, 0, 5, 5, 5, 0, 0, 5, 5, 5, 5, 3, 0, 0, 0, 3, 0, 0 }, 
'{ 0, 0, 0, 3, 3, 5, 5, 5, 0, 5, 5, 5, 5, 5, 5, 0, 5, 0, 5, 5, 0, 5, 5, 0, 0, 3, 3, 0, 0, 0, 3, 3 }, 
'{ 0, 0, 0, 3, 3, 5, 5, 5, 5, 0, 5, 5, 6, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 0, 3, 3, 3, 3, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 3, 3, 3, 3, 3, 0, 5, 5, 5, 5, 6, 5, 5, 5, 5, 5, 5, 6, 5, 5, 0, 5, 3, 3, 3, 0, 0, 0 }, 
'{ 0, 0, 6, 0, 0, 3, 3, 3, 3, 3, 0, 5, 0, 5, 5, 0, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 3, 3, 0, 0, 0 }, 
'{ 0, 3, 0, 0, 0, 0, 0, 3, 3, 3, 0, 5, 5, 0, 0, 5, 5, 5, 5, 0, 5, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 6, 0, 0, 3, 3, 0, 3, 3, 3, 5, 5, 5, 5, 5, 5, 5, 3, 3, 0, 3, 3, 3, 3, 0, 0, 5, 5, 0 }, 
'{ 0, 0, 0, 3, 3, 3, 0, 0, 0, 0, 3, 3, 3, 3, 3, 3, 5, 0, 5, 5, 3, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0 }, 
'{ 0, 0, 6, 6, 0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 3, 5, 5, 5, 3, 3, 0, 0, 0, 0, 0, 6, 0, 6, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0 }, 
'{ 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3 } 
};

explosion_3 <= 
'{ 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 5, 0, 0, 0 }, 
'{ 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 5, 5, 0, 6, 5, 3, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 5, 5, 0, 0, 0, 0, 5, 3, 3, 5, 5, 5, 5, 5, 0, 0, 0, 3, 0, 0, 0, 6, 5, 5, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 5, 0, 5, 0, 0, 5, 5, 5, 3, 0, 5, 0, 5, 5, 0, 0, 0, 5, 5, 0, 6, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 5, 0, 0, 5, 5, 0, 5, 0, 5, 0, 3, 3, 5, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 5, 5, 0, 0, 0, 5, 5, 5, 0, 5, 6, 3, 3, 3, 3, 5, 5, 5, 0, 0, 5, 5, 5, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 5, 0, 5, 5, 5, 5, 5, 0, 5, 5, 0, 3, 5, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 5, 0, 0, 0, 3, 5, 5, 0, 5, 6, 5, 5, 5, 5, 5, 5, 5, 3, 5, 3, 5, 3, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 3, 3, 0, 0, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 6, 5, 0, 5, 3, 0, 0, 5, 5, 5, 0, 0, 0 }, 
'{ 0, 0, 0, 5, 5, 5, 0, 5, 0, 5, 5, 0, 0, 5, 5, 5, 5, 0, 5, 6, 5, 5, 0, 5, 3, 0, 0, 5, 0, 0, 0, 0 }, 
'{ 0, 0, 3, 5, 5, 0, 5, 5, 5, 0, 5, 0, 5, 0, 5, 0, 0, 5, 5, 5, 5, 5, 0, 5, 5, 0, 0, 6, 5, 0, 0, 0 }, 
'{ 0, 0, 3, 5, 0, 5, 5, 5, 5, 5, 5, 5, 0, 5, 0, 5, 0, 5, 5, 5, 5, 0, 5, 5, 5, 0, 6, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 5, 3, 0, 5, 5, 5, 0, 5, 5, 5, 0, 0, 5, 6, 0, 0, 0, 5, 5, 5, 5, 3, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 6, 5, 0, 5, 5, 5, 0, 0, 0, 0, 5, 5, 5, 5, 5, 5, 0, 0, 5, 5, 3, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 3, 6, 0, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 0, 0, 0, 0, 5, 5, 5, 5, 5, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 3, 5, 5, 0, 5, 5, 5, 5, 5, 0, 0, 0, 5, 5, 5, 0, 5, 5, 5, 5, 0, 3, 5, 3, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 3, 5, 3, 5, 5, 5, 5, 0, 5, 5, 0, 6, 0, 5, 0, 5, 5, 5, 5, 5, 5, 0, 5, 3, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 5, 5, 5, 5, 0, 5, 5, 5, 0, 5, 0, 0, 0, 0, 0, 5, 5, 5, 5, 0, 5, 5, 3, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 5, 3, 5, 5, 0, 5, 5, 0, 0, 0, 5, 5, 0, 5, 5, 0, 5, 6, 5, 5, 0, 3, 5, 0, 6, 0, 0, 0, 0 }, 
'{ 0, 5, 0, 0, 3, 5, 0, 5, 5, 5, 0, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 0, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 5, 0, 0, 0, 3, 5, 5, 5, 5, 5, 3, 3, 5, 5, 5, 5, 5, 5, 5, 0, 3, 5, 3, 0, 3, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 3, 5, 5, 5, 5, 5, 5, 6, 5, 5, 5, 5, 5, 0, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 5, 5, 0, 0, 3, 3, 0, 5, 5, 0, 5, 5, 5, 5, 0, 5, 5, 5, 0, 0, 5, 5, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 5, 0, 0, 5, 0, 0, 3, 5, 0, 0, 3, 3, 0, 5, 5, 5, 0, 5, 3, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 5, 0, 5, 0, 0, 5, 3, 3, 3, 5, 5, 0, 3, 3, 5, 5, 3, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 5, 0, 0, 5, 0, 0, 0, 5, 5, 0, 5, 5, 0, 0, 0, 5, 3, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0 }, 
'{ 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 5, 5, 5, 5, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 5, 5, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 }, 
'{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 } 
};
  
  	
	

end	
endmodule